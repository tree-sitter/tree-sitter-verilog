module add ();

endmodule
